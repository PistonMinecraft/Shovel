module constant

pub interface RefInfo {
	class_index u16
	name_and_type_index u16
}
