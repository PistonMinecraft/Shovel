module annotation

pub enum PrimitiveType {
	boolean
	byte
	char
	double
	float
	int
	long
	short
}
