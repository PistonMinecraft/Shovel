module modules

import shovel.reader.constant

pub fn read_module_packages(info []u8, pool constant.ConstantPool) ?[]constant.ConstantPackageInfo {
	return none // TODO
}

pub fn read_module_main_class(info []u8, pool constant.ConstantPool) ?constant.ConstantClassInfo {
	return none // TODO
}
