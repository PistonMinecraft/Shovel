module constant

pub interface DynamicInfo {
	bootstrap_method_attr_index u16
	name_and_type_index         u16
}
